** sch_path: /home/kafkayash/sram_6T_cell/sram_6t_cell.sch
**.subckt sram_6t_cell BL WL BLB Q Qbar
*.ipin BL
*.ipin WL
*.ipin BLB
*.ipin Q
*.opin Qbar
XM26 Q Qbar VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM17 Q Qbar GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM1 Qbar Q GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM2 Qbar Q VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
VDD VDD GND 1.8
XM3 BL WL Q GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM4 BLB WL Qbar GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
vblb BLB GND pulse(1 0 0 10ns 10ns 50ns 100ns)
vbl BL GND pulse(0 1 0 10ns 10ns 50ns 100ns)
vwl WL GND pulse(0 1.3 0 10ns 10ns 50ns 100ns)
Vin Q GND 0
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



 .dc Vin 0 1.8 0.01

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
