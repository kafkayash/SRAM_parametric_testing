* sch_path: /home/yashwanth/sram_6T_cell/sram_6t_cell.sch
**.subckt sram_6t_cell BL WL BLB Q Qbar
*.ipin BL
*.ipin WL
*.ipin BLB
*.ipin Q
*.opin Qbar
XM26 Q Qbar VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L_pmos} W={W_pmos} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 Q Qbar GND GND sky130_fd_pr__nfet_01v8_lvt L={L_nmos} W={W_nmos} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Qbar Q GND GND sky130_fd_pr__nfet_01v8_lvt L={L_nmos} W={W_nmos} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Qbar Q VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L_pmos} W={W_pmos} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VDD VDD GND 1.8
XM3 BL WL Q GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 BLB WL Qbar GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
vblb BLB GND pulse(1 0 0 10ns 10ns 50ns 100ns)
vbl BL GND pulse(0 1 0 10ns 10ns 50ns 100ns)
vwl WL GND pulse(0 1.3 0 10ns 10ns 50ns 100ns)
Vin Q GND 0
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



 .dc Vin 0 1.8 0.01

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
.control
 run
let dVQbar=deriv(V(Qbar))
meas dc Vil FIND V(Q) WHEN dVQbar=-1 CROSS=1
meas dc Vih FIND V(Q) WHEN dVQbar=-1 CROSS=2
meas dc Vol FIND V(Qbar) WHEN dVQbar=-1 CROSS=2
meas dc Voh FIND V(Qbar) AT=0.1
let NM_H=Voh-Vih
let NM_L=Vil-Vol
print NM_L NM_H
.endc                                                                                                                                                                                                        

